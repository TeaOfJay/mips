module cache_decoder(
	input[6:0] addr,
	output reg [127:0] enable
);

always @(addr) begin
	case(addr) 
		7'h01: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0001;
		7'h02: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0002;
		7'h03: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0004;
		7'h04: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0008;
		7'h05: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0010;
		7'h06: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0020;
		7'h07: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0040;
		7'h08: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0080;
		7'h09: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0100;
		7'h0A: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0200;
		7'h0B: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0400;
		7'h0C: enable = 128'h0000_0000_0000_0000_0000_0000_0000_0800;
		7'h0D: enable = 128'h0000_0000_0000_0000_0000_0000_0000_1000;
		7'h0E: enable = 128'h0000_0000_0000_0000_0000_0000_0000_2000;
		7'h0F: enable = 128'h0000_0000_0000_0000_0000_0000_0000_4000;
		7'h10: enable = 128'h0000_0000_0000_0000_0000_0000_0000_8000;
		7'h11: enable = 128'h0000_0000_0000_0000_0000_0000_0001_0000;
		7'h12: enable = 128'h0000_0000_0000_0000_0000_0000_0002_0000;
		7'h13: enable = 128'h0000_0000_0000_0000_0000_0000_0004_0000;
		7'h14: enable = 128'h0000_0000_0000_0000_0000_0000_0008_0000;
		7'h15: enable = 128'h0000_0000_0000_0000_0000_0000_0010_0000;
		7'h16: enable = 128'h0000_0000_0000_0000_0000_0000_0020_0000;
		7'h17: enable = 128'h0000_0000_0000_0000_0000_0000_0040_0000;
		7'h18: enable = 128'h0000_0000_0000_0000_0000_0000_0080_0000;
		7'h19: enable = 128'h0000_0000_0000_0000_0000_0000_0100_0000;
		7'h1A: enable = 128'h0000_0000_0000_0000_0000_0000_0200_0000;
		7'h1B: enable = 128'h0000_0000_0000_0000_0000_0000_0400_0000;
		7'h1C: enable = 128'h0000_0000_0000_0000_0000_0000_0800_0000;
		7'h1D: enable = 128'h0000_0000_0000_0000_0000_0000_1000_0000;
		7'h1E: enable = 128'h0000_0000_0000_0000_0000_0000_2000_0000;
		7'h1F: enable = 128'h0000_0000_0000_0000_0000_0000_4000_0000;
		7'h21: enable = 128'h0000_0000_0000_0000_0000_0000_8000_0000;
		7'h22: enable = 128'h0000_0000_0000_0000_0000_0001_0000_0000;
		7'h23: enable = 128'h0000_0000_0000_0000_0000_0002_0000_0000;
		7'h24: enable = 128'h0000_0000_0000_0000_0000_0004_0000_0000;
		7'h25: enable = 128'h0000_0000_0000_0000_0000_0008_0000_0000;
		7'h26: enable = 128'h0000_0000_0000_0000_0000_0010_0000_0000;
		7'h27: enable = 128'h0000_0000_0000_0000_0000_0020_0000_0000;
		7'h28: enable = 128'h0000_0000_0000_0000_0000_0040_0000_0000;
		7'h29: enable = 128'h0000_0000_0000_0000_0000_0080_0000_0000;
		7'h2A: enable = 128'h0000_0000_0000_0000_0000_0100_0000_0000;
		7'h2B: enable = 128'h0000_0000_0000_0000_0000_0200_0000_0000;
		7'h2C: enable = 128'h0000_0000_0000_0000_0000_0400_0000_0000;
		7'h2D: enable = 128'h0000_0000_0000_0000_0000_0800_0000_0000;
		7'h2E: enable = 128'h0000_0000_0000_0000_0000_1000_0000_0000;
		7'h2F: enable = 128'h0000_0000_0000_0000_0000_2000_0000_0000;
		7'h30: enable = 128'h0000_0000_0000_0000_0000_4000_0000_0000;
		7'h31: enable = 128'h0000_0000_0000_0000_0000_8000_0000_0000;
		7'h32: enable = 128'h0000_0000_0000_0000_0001_0000_0000_0000;
		7'h33: enable = 128'h0000_0000_0000_0000_0002_0000_0000_0000;
		7'h34: enable = 128'h0000_0000_0000_0000_0004_0000_0000_0000;
		7'h35: enable = 128'h0000_0000_0000_0000_0008_0000_0000_0000;
		7'h36: enable = 128'h0000_0000_0000_0000_0010_0000_0000_0000;
		7'h37: enable = 128'h0000_0000_0000_0000_0020_0000_0000_0000;
		7'h38: enable = 128'h0000_0000_0000_0000_0040_0000_0000_0000;
		7'h39: enable = 128'h0000_0000_0000_0000_0080_0000_0000_0000;
		7'h3A: enable = 128'h0000_0000_0000_0000_0100_0000_0000_0000;
		7'h3B: enable = 128'h0000_0000_0000_0000_0200_0000_0000_0000;
		7'h3C: enable = 128'h0000_0000_0000_0000_0400_0000_0000_0000;
		7'h3D: enable = 128'h0000_0000_0000_0000_0800_0000_0000_0000;
		7'h3E: enable = 128'h0000_0000_0000_0000_1000_0000_0000_0000;
		7'h3F: enable = 128'h0000_0000_0000_0000_2000_0000_0000_0000;
		7'h40: enable = 128'h0000_0000_0000_0000_4000_0000_0000_0000;
		7'h41: enable = 128'h0000_0000_0000_0000_8000_0000_0000_0000;
		7'h42: enable = 128'h0000_0000_0000_0001_0000_0000_0000_0000;
		7'h43: enable = 128'h0000_0000_0000_0002_0000_0000_0000_0000;
		7'h44: enable = 128'h0000_0000_0000_0004_0000_0000_0000_0000;
		7'h45: enable = 128'h0000_0000_0000_0008_0000_0000_0000_0000;
		7'h46: enable = 128'h0000_0000_0000_0010_0000_0000_0000_0000;
		7'h47: enable = 128'h0000_0000_0000_0020_0000_0000_0000_0000;
		7'h48: enable = 128'h0000_0000_0000_0040_0000_0000_0000_0000;
		7'h49: enable = 128'h0000_0000_0000_0080_0000_0000_0000_0000;
		7'h4A: enable = 128'h0000_0000_0000_0100_0000_0000_0000_0000;
		7'h4B: enable = 128'h0000_0000_0000_0200_0000_0000_0000_0000;
		7'h4C: enable = 128'h0000_0000_0000_0400_0000_0000_0000_0000;
		7'h4D: enable = 128'h0000_0000_0000_0800_0000_0000_0000_0000;
		7'h4E: enable = 128'h0000_0000_0000_1000_0000_0000_0000_0000;
		7'h4F: enable = 128'h0000_0000_0000_2000_0000_0000_0000_0000;
		7'h50: enable = 128'h0000_0000_0000_4000_0000_0000_0000_0000;
		7'h51: enable = 128'h0000_0000_0000_8000_0000_0000_0000_0000;
		7'h52: enable = 128'h0000_0000_0001_0000_0000_0000_0000_0000;
		7'h53: enable = 128'h0000_0000_0002_0000_0000_0000_0000_0000;
		7'h54: enable = 128'h0000_0000_0004_0000_0000_0000_0000_0000;
		7'h55: enable = 128'h0000_0000_0008_0000_0000_0000_0000_0000;
		7'h56: enable = 128'h0000_0000_0010_0000_0000_0000_0000_0000;
		7'h57: enable = 128'h0000_0000_0020_0000_0000_0000_0000_0000;
		7'h58: enable = 128'h0000_0000_0040_0000_0000_0000_0000_0000;
		7'h59: enable = 128'h0000_0000_0080_0000_0000_0000_0000_0000;
		7'h5A: enable = 128'h0000_0000_0100_0000_0000_0000_0000_0000;
		7'h5B: enable = 128'h0000_0000_0200_0000_0000_0000_0000_0000;
		7'h5C: enable = 128'h0000_0000_0400_0000_0000_0000_0000_0000;
		7'h5D: enable = 128'h0000_0000_0800_0000_0000_0000_0000_0000;
		7'h5E: enable = 128'h0000_0000_1000_0000_0000_0000_0000_0000;
		7'h5F: enable = 128'h0000_0000_2000_0000_0000_0000_0000_0000;
		7'h60: enable = 128'h0000_0000_4000_0000_0000_0000_0000_0000;
		7'h61: enable = 128'h0000_0000_8000_0000_0000_0000_0000_0000;
		7'h62: enable = 128'h0000_0001_0000_0000_0000_0000_0000_0000;
		7'h63: enable = 128'h0000_0002_0000_0000_0000_0000_0000_0000;
		7'h64: enable = 128'h0000_0004_0000_0000_0000_0000_0000_0000;
		7'h65: enable = 128'h0000_0008_0000_0000_0000_0000_0000_0000;
		7'h66: enable = 128'h0000_0010_0000_0000_0000_0000_0000_0000;
		7'h67: enable = 128'h0000_0020_0000_0000_0000_0000_0000_0000;
		7'h68: enable = 128'h0000_0040_0000_0000_0000_0000_0000_0000;
		7'h69: enable = 128'h0000_0080_0000_0000_0000_0000_0000_0000;
		7'h6A: enable = 128'h0000_0100_0000_0000_0000_0000_0000_0000;
		7'h6B: enable = 128'h0000_0200_0000_0000_0000_0000_0000_0000;
		7'h6C: enable = 128'h0000_0400_0000_0000_0000_0000_0000_0000;
		7'h6D: enable = 128'h0000_0800_0000_0000_0000_0000_0000_0000;
		7'h6E: enable = 128'h0000_1000_0000_0000_0000_0000_0000_0000;
		7'h6F: enable = 128'h0000_2000_0000_0000_0000_0000_0000_0000;
		7'h70: enable = 128'h0000_4000_0000_0000_0000_0000_0000_0000;
		7'h71: enable = 128'h0000_8000_0000_0000_0000_0000_0000_0000;
		7'h72: enable = 128'h0001_0000_0000_0000_0000_0000_0000_0000;
		7'h73: enable = 128'h0002_0000_0000_0000_0000_0000_0000_0000;
		7'h74: enable = 128'h0004_0000_0000_0000_0000_0000_0000_0000;
		7'h75: enable = 128'h0008_0000_0000_0000_0000_0000_0000_0000;
		7'h76: enable = 128'h0010_0000_0000_0000_0000_0000_0000_0000;
		7'h77: enable = 128'h0020_0000_0000_0000_0000_0000_0000_0000;
		7'h78: enable = 128'h0040_0000_0000_0000_0000_0000_0000_0000;
		7'h79: enable = 128'h0080_0000_0000_0000_0000_0000_0000_0000;
		7'h7A: enable = 128'h0100_0000_0000_0000_0000_0000_0000_0000;
		7'h7B: enable = 128'h0200_0000_0000_0000_0000_0000_0000_0000;
		7'h7C: enable = 128'h0400_0000_0000_0000_0000_0000_0000_0000;
		7'h7D: enable = 128'h0800_0000_0000_0000_0000_0000_0000_0000;
		7'h7E: enable = 128'h1000_0000_0000_0000_0000_0000_0000_0000;
		7'h7F: enable = 128'h2000_0000_0000_0000_0000_0000_0000_0000;
		default: enable = 128'h0;
	endcase // addr
end

endmodule // cache_decoder