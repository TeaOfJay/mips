module idex(

input[15:0] q_reg1,
input[15:0] q_reg2,


output[15:0] d_reg1,
output[15:0] d_reg2
	);



endmodule // idex